library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity example is
    port (

    );
end entity example;

architecture bhv of example is
begin

end bhv;